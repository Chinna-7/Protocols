interface 


endinterface
