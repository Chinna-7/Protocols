`include "spi_interface.sv"
`include "spi_seq_item.sv"
`include "spi_seq.sv"
`include "spi_seqr.sv"
`include "spi_driver.sv"
`include "spi_monitor.sv"
`include "spi_agent.sv"
`include "spi_scoreboard1.sv"
`include "spi_scoreboard2.sv"
`include "spi_environment.sv"
`include "spi_test.sv"